library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
-- using " word address " below
-- system instruction area : 0x0000 ~ 0x3fff
-- user instruction area : 0x4000 ~ 0x7fff
-- system data area : 0x8000 ~ 0xbeff
-- com1 : 0xbf00 ~ 0xbf01
-- com2 : 0xbf02 ~ 0xbf03
-- resident : 0xbf04 ~ 0xbf0f
-- system heap stack : 0xbf10 ~ 0xbfff
-- user data area : 0xc000 ~ 0xffff
entity memory is
	port(
		LFlag, SFlag : in std_logic;
		Address : in std_logic_vector(15 downto 0);
		DataS : in std_logic_vector(15 downto 0);
		InstructionAddress : in std_logic_vector(15 downto 0);
		clk : in std_logic;
		clk_scan : in std_logic;
		reset : in std_logic;
		
		Result : out std_logic_vector(15 downto 0);
        Result_L_pointer : out std_logic;
        Result_L : out std_logic_vector(15 downto 0);
		InstructionResult : out std_logic_vector(15 downto 0);

		-- data mem
		Ram1Data : inout std_logic_vector(15 downto 0);
		Ram1Addr : out std_logic_vector(15 downto 0);
		Ram1OE, Ram1WE, Ram1EN : out std_logic;
		dataReady, rdn, wrn, tbre, tsre : inout std_logic;

		-- instruction mem
		Ram2Data : inout std_logic_vector(15 downto 0);
		Ram2Addr : out std_logic_vector(15 downto 0);
		Ram2OE, Ram2WE, Ram2EN : out std_logic;
		
		-- flash
		flashByte : out std_logic;
		flashVpen : out std_logic;
		flashCE : out std_logic;
		flashOE : out std_logic;
		flashWE : out std_logic;
		flashRP : out std_logic;
		flashAddr : out std_logic_vector(22 downto 1);
		flashData : inout std_logic_vector(15 downto 0);
		
		-- led
		led : out std_logic_vector(15 downto 0);
		started : out std_logic
		--trigger : out std_logic_vector(49 downto 0)
	);
end memory;

architecture bhv of memory is
type ramBlock is array(1023 downto 0) of std_logic_vector(15 downto 0);
signal Ram1, Ram2 : ramBlock;

-- instruction [0000,0013]
-- data [c000,c013]
signal startedCache : std_logic := '0';
signal triggerCache : std_logic_vector(49 downto 0) := (others => '1');
begin
	started <= startedCache;
	--trigger <= triggerCache;
	led <= (others => '0');
	process (LFlag, SFlag, startedCache, clk_scan, clk, reset)
	begin
		if (reset = '1') then
			startedCache <= '1';
            Ram2(0) <= x"1002";
            Ram2(1) <= x"0800";
            Ram2(2) <= x"0800";
            Ram2(3) <= x"1002";
            Ram2(4) <= x"0800";
            Ram2(5) <= x"0800";
            Ram2(6) <= x"ef40";
            Ram2(7) <= x"4f03";
            Ram2(8) <= x"0000";
            Ram2(9) <= x"0000";
            Ram2(10) <= x"0000";
            Ram2(11) <= x"0000";
            Ram2(12) <= x"0000";
            Ram2(13) <= x"0000";
            Ram2(14) <= x"0000";
            Ram2(15) <= x"0000";
            Ram2(16) <= x"0000";
            Ram2(17) <= x"0000";
            Ram2(18) <= x"0000";
            Ram2(19) <= x"0000";
            Ram2(20) <= x"0000";
            Ram2(21) <= x"0000";
            Ram2(22) <= x"0000";
            Ram2(23) <= x"0000";
            Ram2(24) <= x"0000";
            Ram2(25) <= x"0000";
            Ram2(26) <= x"0000";
            Ram2(27) <= x"0000";
            Ram2(28) <= x"0000";
            Ram2(29) <= x"0000";
            Ram2(30) <= x"0000";
            Ram2(31) <= x"0000";
            Ram2(32) <= x"0000";
            Ram2(33) <= x"0000";
            Ram2(34) <= x"0000";
            Ram2(35) <= x"0000";
            Ram2(36) <= x"0000";
            Ram2(37) <= x"0000";
            Ram2(38) <= x"0000";
            Ram2(39) <= x"0000";
            Ram2(40) <= x"0000";
            Ram2(41) <= x"0000";
            Ram2(42) <= x"0000";
            Ram2(43) <= x"0000";
            Ram2(44) <= x"0000";
            Ram2(45) <= x"0000";
            Ram2(46) <= x"0000";
            Ram2(47) <= x"0000";
            Ram2(48) <= x"0000";
            Ram2(49) <= x"0000";
            Ram2(50) <= x"0000";
            Ram2(51) <= x"0000";
            Ram2(52) <= x"0000";
            Ram2(53) <= x"0000";
            Ram2(54) <= x"0000";
            Ram2(55) <= x"0000";
            Ram2(56) <= x"0000";
            Ram2(57) <= x"0000";
            Ram2(58) <= x"0000";
            Ram2(59) <= x"0000";
            Ram2(60) <= x"0000";
            Ram2(61) <= x"0000";
            Ram2(62) <= x"0000";
            Ram2(63) <= x"0000";
            Ram2(64) <= x"0000";
            Ram2(65) <= x"0000";
            Ram2(66) <= x"0000";
            Ram2(67) <= x"0000";
            Ram2(68) <= x"0000";
            Ram2(69) <= x"0000";
            Ram2(70) <= x"0000";
            Ram2(71) <= x"0000";
            Ram2(72) <= x"0000";
            Ram2(73) <= x"0000";
            Ram2(74) <= x"0000";
            Ram2(75) <= x"0000";
            Ram2(76) <= x"0000";
            Ram2(77) <= x"0000";
            Ram2(78) <= x"0000";
            Ram2(79) <= x"0000";
            Ram2(80) <= x"0000";
            Ram2(81) <= x"0000";
            Ram2(82) <= x"0000";
            Ram2(83) <= x"0000";
            Ram2(84) <= x"0000";
            Ram2(85) <= x"0000";
            Ram2(86) <= x"0000";
            Ram2(87) <= x"0000";
            Ram2(88) <= x"0000";
            Ram2(89) <= x"0000";
            Ram2(90) <= x"0000";
            Ram2(91) <= x"0000";
            Ram2(92) <= x"0000";
            Ram2(93) <= x"0000";
            Ram2(94) <= x"0000";
            Ram2(95) <= x"0000";
            Ram2(96) <= x"0000";
            Ram2(97) <= x"0000";
            Ram2(98) <= x"0000";
            Ram2(99) <= x"0000";
            Ram2(100) <= x"0000";
            Ram2(101) <= x"0000";
            Ram2(102) <= x"0000";
            Ram2(103) <= x"0000";
            Ram2(104) <= x"0000";
            Ram2(105) <= x"0000";
            Ram2(106) <= x"0000";
            Ram2(107) <= x"0000";
            Ram2(108) <= x"0000";
            Ram2(109) <= x"0000";
            Ram2(110) <= x"0000";
            Ram2(111) <= x"0000";
            Ram2(112) <= x"0000";
            Ram2(113) <= x"0000";
            Ram2(114) <= x"0000";
            Ram2(115) <= x"0000";
            Ram2(116) <= x"0000";
            Ram2(117) <= x"0000";
            Ram2(118) <= x"0000";
            Ram2(119) <= x"0000";
            Ram2(120) <= x"0000";
            Ram2(121) <= x"0000";
            Ram2(122) <= x"0000";
            Ram2(123) <= x"0000";
            Ram2(124) <= x"0000";
            Ram2(125) <= x"0000";
            Ram2(126) <= x"0000";
            Ram2(127) <= x"0000";
            Ram2(128) <= x"0000";
            Ram2(129) <= x"0000";
            Ram2(130) <= x"0000";
            Ram2(131) <= x"0000";
            Ram2(132) <= x"0000";
            Ram2(133) <= x"0000";
            Ram2(134) <= x"0000";
            Ram2(135) <= x"0000";
            Ram2(136) <= x"0000";
            Ram2(137) <= x"0000";
            Ram2(138) <= x"0000";
            Ram2(139) <= x"0000";
            Ram2(140) <= x"0000";
            Ram2(141) <= x"0000";
            Ram2(142) <= x"0000";
            Ram2(143) <= x"0000";
            Ram2(144) <= x"0000";
            Ram2(145) <= x"0000";
            Ram2(146) <= x"0000";
            Ram2(147) <= x"0000";
            Ram2(148) <= x"0000";
            Ram2(149) <= x"0000";
            Ram2(150) <= x"0000";
            Ram2(151) <= x"0000";
            Ram2(152) <= x"0000";
            Ram2(153) <= x"0000";
            Ram2(154) <= x"0000";
            Ram2(155) <= x"0000";
            Ram2(156) <= x"0000";
            Ram2(157) <= x"0000";
            Ram2(158) <= x"0000";
            Ram2(159) <= x"0000";
            Ram2(160) <= x"0000";
            Ram2(161) <= x"0000";
            Ram2(162) <= x"0000";
            Ram2(163) <= x"0000";
            Ram2(164) <= x"0000";
            Ram2(165) <= x"0000";
            Ram2(166) <= x"0000";
            Ram2(167) <= x"0000";
            Ram2(168) <= x"0000";
            Ram2(169) <= x"0000";
            Ram2(170) <= x"0000";
            Ram2(171) <= x"0000";
            Ram2(172) <= x"0000";
            Ram2(173) <= x"0000";
            Ram2(174) <= x"0000";
            Ram2(175) <= x"0000";
            Ram2(176) <= x"0000";
            Ram2(177) <= x"0000";
            Ram2(178) <= x"0000";
            Ram2(179) <= x"0000";
            Ram2(180) <= x"0000";
            Ram2(181) <= x"0000";
            Ram2(182) <= x"0000";
            Ram2(183) <= x"0000";
            Ram2(184) <= x"0000";
            Ram2(185) <= x"0000";
            Ram2(186) <= x"0000";
            Ram2(187) <= x"0000";
            Ram2(188) <= x"0000";
            Ram2(189) <= x"0000";
            Ram2(190) <= x"0000";
            Ram2(191) <= x"0000";
            Ram2(192) <= x"0000";
            Ram2(193) <= x"0000";
            Ram2(194) <= x"0000";
            Ram2(195) <= x"0000";
            Ram2(196) <= x"0000";
            Ram2(197) <= x"0000";
            Ram2(198) <= x"0000";
            Ram2(199) <= x"0000";
            Ram2(200) <= x"0000";
            Ram2(201) <= x"0000";
            Ram2(202) <= x"0000";
            Ram2(203) <= x"0000";
            Ram2(204) <= x"0000";
            Ram2(205) <= x"0000";
            Ram2(206) <= x"0000";
            Ram2(207) <= x"0000";
            Ram2(208) <= x"0000";
            Ram2(209) <= x"0000";
            Ram2(210) <= x"0000";
            Ram2(211) <= x"0000";
            Ram2(212) <= x"0000";
            Ram2(213) <= x"0000";
            Ram2(214) <= x"0000";
            Ram2(215) <= x"0000";
            Ram2(216) <= x"0000";
            Ram2(217) <= x"0000";
            Ram2(218) <= x"0000";
            Ram2(219) <= x"0000";
            Ram2(220) <= x"0000";
            Ram2(221) <= x"0000";
            Ram2(222) <= x"0000";
            Ram2(223) <= x"0000";
            Ram2(224) <= x"0000";
            Ram2(225) <= x"0000";
            Ram2(226) <= x"0000";
            Ram2(227) <= x"0000";
            Ram2(228) <= x"0000";
            Ram2(229) <= x"0000";
            Ram2(230) <= x"0000";
            Ram2(231) <= x"0000";
            Ram2(232) <= x"0000";
            Ram2(233) <= x"0000";
            Ram2(234) <= x"0000";
            Ram2(235) <= x"0000";
            Ram2(236) <= x"0000";
            Ram2(237) <= x"0000";
            Ram2(238) <= x"0000";
            Ram2(239) <= x"0000";
            Ram2(240) <= x"0000";
            Ram2(241) <= x"0000";
            Ram2(242) <= x"0000";
            Ram2(243) <= x"0000";
            Ram2(244) <= x"0000";
            Ram2(245) <= x"0000";
            Ram2(246) <= x"0000";
            Ram2(247) <= x"0000";
            Ram2(248) <= x"0000";
            Ram2(249) <= x"0000";
            Ram2(250) <= x"0000";
            Ram2(251) <= x"0000";
            Ram2(252) <= x"0000";
            Ram2(253) <= x"0000";
            Ram2(254) <= x"0000";
            Ram2(255) <= x"0000";
            Ram2(256) <= x"0000";
            Ram2(257) <= x"0000";
            Ram2(258) <= x"0000";
            Ram2(259) <= x"0000";
            Ram2(260) <= x"0000";
            Ram2(261) <= x"0000";
            Ram2(262) <= x"0000";
            Ram2(263) <= x"0000";
            Ram2(264) <= x"0000";
            Ram2(265) <= x"0000";
            Ram2(266) <= x"0000";
            Ram2(267) <= x"0000";
            Ram2(268) <= x"0000";
            Ram2(269) <= x"0000";
            Ram2(270) <= x"0000";
            Ram2(271) <= x"0000";
            Ram2(272) <= x"0000";
            Ram2(273) <= x"0000";
            Ram2(274) <= x"0000";
            Ram2(275) <= x"0000";
            Ram2(276) <= x"0000";
            Ram2(277) <= x"0000";
            Ram2(278) <= x"0000";
            Ram2(279) <= x"0000";
            Ram2(280) <= x"0000";
            Ram2(281) <= x"0000";
            Ram2(282) <= x"0000";
            Ram2(283) <= x"0000";
            Ram2(284) <= x"0000";
            Ram2(285) <= x"0000";
            Ram2(286) <= x"0000";
            Ram2(287) <= x"0000";
            Ram2(288) <= x"0000";
            Ram2(289) <= x"0000";
            Ram2(290) <= x"0000";
            Ram2(291) <= x"0000";
            Ram2(292) <= x"0000";
            Ram2(293) <= x"0000";
            Ram2(294) <= x"0000";
            Ram2(295) <= x"0000";
            Ram2(296) <= x"0000";
            Ram2(297) <= x"0000";
            Ram2(298) <= x"0000";
            Ram2(299) <= x"0000";
            Ram2(300) <= x"0000";
            Ram2(301) <= x"0000";
            Ram2(302) <= x"0000";
            Ram2(303) <= x"0000";
            Ram2(304) <= x"0000";
            Ram2(305) <= x"0000";
            Ram2(306) <= x"0000";
            Ram2(307) <= x"0000";
            Ram2(308) <= x"0000";
            Ram2(309) <= x"0000";
            Ram2(310) <= x"0000";
            Ram2(311) <= x"0000";
            Ram2(312) <= x"0000";
            Ram2(313) <= x"0000";
            Ram2(314) <= x"0000";
            Ram2(315) <= x"0000";
            Ram2(316) <= x"0000";
            Ram2(317) <= x"0000";
            Ram2(318) <= x"0000";
            Ram2(319) <= x"0000";
            Ram2(320) <= x"0000";
            Ram2(321) <= x"0000";
            Ram2(322) <= x"0000";
            Ram2(323) <= x"0000";
            Ram2(324) <= x"0000";
            Ram2(325) <= x"0000";
            Ram2(326) <= x"0000";
            Ram2(327) <= x"0000";
            Ram2(328) <= x"0000";
            Ram2(329) <= x"0000";
            Ram2(330) <= x"0000";
            Ram2(331) <= x"0000";
            Ram2(332) <= x"0000";
            Ram2(333) <= x"0000";
            Ram2(334) <= x"0000";
            Ram2(335) <= x"0000";
            Ram2(336) <= x"0000";
            Ram2(337) <= x"0000";
            Ram2(338) <= x"0000";
            Ram2(339) <= x"0000";
            Ram2(340) <= x"0000";
            Ram2(341) <= x"0000";
            Ram2(342) <= x"0000";
            Ram2(343) <= x"0000";
            Ram2(344) <= x"0000";
            Ram2(345) <= x"0000";
            Ram2(346) <= x"0000";
            Ram2(347) <= x"0000";
            Ram2(348) <= x"0000";
            Ram2(349) <= x"0000";
            Ram2(350) <= x"0000";
            Ram2(351) <= x"0000";
            Ram2(352) <= x"0000";
            Ram2(353) <= x"0000";
            Ram2(354) <= x"0000";
            Ram2(355) <= x"0000";
            Ram2(356) <= x"0000";
            Ram2(357) <= x"0000";
            Ram2(358) <= x"0000";
            Ram2(359) <= x"0000";
            Ram2(360) <= x"0000";
            Ram2(361) <= x"0000";
            Ram2(362) <= x"0000";
            Ram2(363) <= x"0000";
            Ram2(364) <= x"0000";
            Ram2(365) <= x"0000";
            Ram2(366) <= x"0000";
            Ram2(367) <= x"0000";
            Ram2(368) <= x"0000";
            Ram2(369) <= x"0000";
            Ram2(370) <= x"0000";
            Ram2(371) <= x"0000";
            Ram2(372) <= x"0000";
            Ram2(373) <= x"0000";
            Ram2(374) <= x"0000";
            Ram2(375) <= x"0000";
            Ram2(376) <= x"0000";
            Ram2(377) <= x"0000";
            Ram2(378) <= x"0000";
            Ram2(379) <= x"0000";
            Ram2(380) <= x"0000";
            Ram2(381) <= x"0000";
            Ram2(382) <= x"0000";
            Ram2(383) <= x"0000";
            Ram2(384) <= x"0000";
            Ram2(385) <= x"0000";
            Ram2(386) <= x"0000";
            Ram2(387) <= x"0000";
            Ram2(388) <= x"0000";
            Ram2(389) <= x"0000";
            Ram2(390) <= x"0000";
            Ram2(391) <= x"0000";
            Ram2(392) <= x"0000";
            Ram2(393) <= x"0000";
            Ram2(394) <= x"0000";
            Ram2(395) <= x"0000";
            Ram2(396) <= x"0000";
            Ram2(397) <= x"0000";
            Ram2(398) <= x"0000";
            Ram2(399) <= x"0000";
            Ram2(400) <= x"0000";
            Ram2(401) <= x"0000";
            Ram2(402) <= x"0000";
            Ram2(403) <= x"0000";
            Ram2(404) <= x"0000";
            Ram2(405) <= x"0000";
            Ram2(406) <= x"0000";
            Ram2(407) <= x"0000";
            Ram2(408) <= x"0000";
            Ram2(409) <= x"0000";
            Ram2(410) <= x"0000";
            Ram2(411) <= x"0000";
            Ram2(412) <= x"0000";
            Ram2(413) <= x"0000";
            Ram2(414) <= x"0000";
            Ram2(415) <= x"0000";
            Ram2(416) <= x"0000";
            Ram2(417) <= x"0000";
            Ram2(418) <= x"0000";
            Ram2(419) <= x"0000";
            Ram2(420) <= x"0000";
            Ram2(421) <= x"0000";
            Ram2(422) <= x"0000";
            Ram2(423) <= x"0000";
            Ram2(424) <= x"0000";
            Ram2(425) <= x"0000";
            Ram2(426) <= x"0000";
            Ram2(427) <= x"0000";
            Ram2(428) <= x"0000";
            Ram2(429) <= x"0000";
            Ram2(430) <= x"0000";
            Ram2(431) <= x"0000";
            Ram2(432) <= x"0000";
            Ram2(433) <= x"0000";
            Ram2(434) <= x"0000";
            Ram2(435) <= x"0000";
            Ram2(436) <= x"0000";
            Ram2(437) <= x"0000";
            Ram2(438) <= x"0000";
            Ram2(439) <= x"0000";
            Ram2(440) <= x"0000";
            Ram2(441) <= x"0000";
            Ram2(442) <= x"0000";
            Ram2(443) <= x"0000";
            Ram2(444) <= x"0000";
            Ram2(445) <= x"0000";
            Ram2(446) <= x"0000";
            Ram2(447) <= x"0000";
            Ram2(448) <= x"0000";
            Ram2(449) <= x"0000";
            Ram2(450) <= x"0000";
            Ram2(451) <= x"0000";
            Ram2(452) <= x"0000";
            Ram2(453) <= x"0000";
            Ram2(454) <= x"0000";
            Ram2(455) <= x"0000";
            Ram2(456) <= x"0000";
            Ram2(457) <= x"0000";
            Ram2(458) <= x"0000";
            Ram2(459) <= x"0000";
            Ram2(460) <= x"0000";
            Ram2(461) <= x"0000";
            Ram2(462) <= x"0000";
            Ram2(463) <= x"0000";
            Ram2(464) <= x"0000";
            Ram2(465) <= x"0000";
            Ram2(466) <= x"0000";
            Ram2(467) <= x"0000";
            Ram2(468) <= x"0000";
            Ram2(469) <= x"0000";
            Ram2(470) <= x"0000";
            Ram2(471) <= x"0000";
            Ram2(472) <= x"0000";
            Ram2(473) <= x"0000";
            Ram2(474) <= x"0000";
            Ram2(475) <= x"0000";
            Ram2(476) <= x"0000";
            Ram2(477) <= x"0000";
            Ram2(478) <= x"0000";
            Ram2(479) <= x"0000";
            Ram2(480) <= x"0000";
            Ram2(481) <= x"0000";
            Ram2(482) <= x"0000";
            Ram2(483) <= x"0000";
            Ram2(484) <= x"0000";
            Ram2(485) <= x"0000";
            Ram2(486) <= x"0000";
            Ram2(487) <= x"0000";
            Ram2(488) <= x"0000";
            Ram2(489) <= x"0000";
            Ram2(490) <= x"0000";
            Ram2(491) <= x"0000";
            Ram2(492) <= x"0000";
            Ram2(493) <= x"0000";
            Ram2(494) <= x"0000";
            Ram2(495) <= x"0000";
            Ram2(496) <= x"0000";
            Ram2(497) <= x"0000";
            Ram2(498) <= x"0000";
            Ram2(499) <= x"0000";
            Ram2(500) <= x"0000";
            Ram2(501) <= x"0000";
            Ram2(502) <= x"0000";
            Ram2(503) <= x"0000";
            Ram2(504) <= x"0000";
            Ram2(505) <= x"0000";
            Ram2(506) <= x"0000";
            Ram2(507) <= x"0000";
            Ram2(508) <= x"0000";
            Ram2(509) <= x"0000";
            Ram2(510) <= x"0000";
            Ram2(511) <= x"0000";
            Ram2(512) <= x"0000";
            Ram2(513) <= x"0000";
            Ram2(514) <= x"0000";
            Ram2(515) <= x"0000";
            Ram2(516) <= x"0000";
            Ram2(517) <= x"0000";
            Ram2(518) <= x"0000";
            Ram2(519) <= x"0000";
            Ram2(520) <= x"0000";
            Ram2(521) <= x"0000";
            Ram2(522) <= x"0000";
            Ram2(523) <= x"0000";
            Ram2(524) <= x"0000";
            Ram2(525) <= x"0000";
            Ram2(526) <= x"0000";
            Ram2(527) <= x"0000";
            Ram2(528) <= x"0000";
            Ram2(529) <= x"0000";
            Ram2(530) <= x"0000";
            Ram2(531) <= x"0000";
            Ram2(532) <= x"0000";
            Ram2(533) <= x"0000";
            Ram2(534) <= x"0000";
            Ram2(535) <= x"0000";
            Ram2(536) <= x"0000";
            Ram2(537) <= x"0000";
            Ram2(538) <= x"0000";
            Ram2(539) <= x"0000";
            Ram2(540) <= x"0000";
            Ram2(541) <= x"0000";
            Ram2(542) <= x"0000";
            Ram2(543) <= x"0000";
            Ram2(544) <= x"0000";
            Ram2(545) <= x"0000";
            Ram2(546) <= x"0000";
            Ram2(547) <= x"0000";
            Ram2(548) <= x"0000";
            Ram2(549) <= x"0000";
            Ram2(550) <= x"0000";
            Ram2(551) <= x"0000";
            Ram2(552) <= x"0000";
            Ram2(553) <= x"0000";
            Ram2(554) <= x"0000";
            Ram2(555) <= x"0000";
            Ram2(556) <= x"0000";
            Ram2(557) <= x"0000";
            Ram2(558) <= x"0000";
            Ram2(559) <= x"0000";
            Ram2(560) <= x"0000";
            Ram2(561) <= x"0000";
            Ram2(562) <= x"0000";
            Ram2(563) <= x"0000";
            Ram2(564) <= x"0000";
            Ram2(565) <= x"0000";
            Ram2(566) <= x"0000";
            Ram2(567) <= x"0000";
            Ram2(568) <= x"0000";
            Ram2(569) <= x"0000";
            Ram2(570) <= x"0000";
            Ram2(571) <= x"0000";
            Ram2(572) <= x"0000";
            Ram2(573) <= x"0000";
            Ram2(574) <= x"0000";
            Ram2(575) <= x"0000";
            Ram2(576) <= x"0000";
            Ram2(577) <= x"0000";
            Ram2(578) <= x"0000";
            Ram2(579) <= x"0000";
            Ram2(580) <= x"0000";
            Ram2(581) <= x"0000";
            Ram2(582) <= x"0000";
            Ram2(583) <= x"0000";
            Ram2(584) <= x"0000";
            Ram2(585) <= x"0000";
            Ram2(586) <= x"0000";
            Ram2(587) <= x"0000";
            Ram2(588) <= x"0000";
            Ram2(589) <= x"0000";
            Ram2(590) <= x"0000";
            Ram2(591) <= x"0000";
            Ram2(592) <= x"0000";
            Ram2(593) <= x"0000";
            Ram2(594) <= x"0000";
            Ram2(595) <= x"0000";
            Ram2(596) <= x"0000";
            Ram2(597) <= x"0000";
            Ram2(598) <= x"0000";
            Ram2(599) <= x"0000";
            Ram2(600) <= x"0000";
            Ram2(601) <= x"0000";
            Ram2(602) <= x"0000";
            Ram2(603) <= x"0000";
            Ram2(604) <= x"0000";
            Ram2(605) <= x"0000";
            Ram2(606) <= x"0000";
            Ram2(607) <= x"0000";
            Ram2(608) <= x"0000";
            Ram2(609) <= x"0000";
            Ram2(610) <= x"0000";
            Ram2(611) <= x"0000";
            Ram2(612) <= x"0000";
            Ram2(613) <= x"0000";
            Ram2(614) <= x"0000";
            Ram2(615) <= x"0000";
            Ram2(616) <= x"0000";
            Ram2(617) <= x"0000";
            Ram2(618) <= x"0000";
            Ram2(619) <= x"0000";
            Ram2(620) <= x"0000";
            Ram2(621) <= x"0000";
            Ram2(622) <= x"0000";
            Ram2(623) <= x"0000";
            Ram2(624) <= x"0000";
            Ram2(625) <= x"0000";
            Ram2(626) <= x"0000";
            Ram2(627) <= x"0000";
            Ram2(628) <= x"0000";
            Ram2(629) <= x"0000";
            Ram2(630) <= x"0000";
            Ram2(631) <= x"0000";
            Ram2(632) <= x"0000";
            Ram2(633) <= x"0000";
            Ram2(634) <= x"0000";
            Ram2(635) <= x"0000";
            Ram2(636) <= x"0000";
            Ram2(637) <= x"0000";
            Ram2(638) <= x"0000";
            Ram2(639) <= x"0000";
            Ram2(640) <= x"0000";
            Ram2(641) <= x"0000";
            Ram2(642) <= x"0000";
            Ram2(643) <= x"0000";
            Ram2(644) <= x"0000";
            Ram2(645) <= x"0000";
            Ram2(646) <= x"0000";
            Ram2(647) <= x"0000";
            Ram2(648) <= x"0000";
            Ram2(649) <= x"0000";
            Ram2(650) <= x"0000";
            Ram2(651) <= x"0000";
            Ram2(652) <= x"0000";
            Ram2(653) <= x"0000";
            Ram2(654) <= x"0000";
            Ram2(655) <= x"0000";
            Ram2(656) <= x"0000";
            Ram2(657) <= x"0000";
            Ram2(658) <= x"0000";
            Ram2(659) <= x"0000";
            Ram2(660) <= x"0000";
            Ram2(661) <= x"0000";
            Ram2(662) <= x"0000";
            Ram2(663) <= x"0000";
            Ram2(664) <= x"0000";
            Ram2(665) <= x"0000";
            Ram2(666) <= x"0000";
            Ram2(667) <= x"0000";
            Ram2(668) <= x"0000";
            Ram2(669) <= x"0000";
            Ram2(670) <= x"0000";
            Ram2(671) <= x"0000";
            Ram2(672) <= x"0000";
            Ram2(673) <= x"0000";
            Ram2(674) <= x"0000";
            Ram2(675) <= x"0000";
            Ram2(676) <= x"0000";
            Ram2(677) <= x"0000";
            Ram2(678) <= x"0000";
            Ram2(679) <= x"0000";
            Ram2(680) <= x"0000";
            Ram2(681) <= x"0000";
            Ram2(682) <= x"0000";
            Ram2(683) <= x"0000";
            Ram2(684) <= x"0000";
            Ram2(685) <= x"0000";
            Ram2(686) <= x"0000";
            Ram2(687) <= x"0000";
            Ram2(688) <= x"0000";
            Ram2(689) <= x"0000";
            Ram2(690) <= x"0000";
            Ram2(691) <= x"0000";
            Ram2(692) <= x"0000";
            Ram2(693) <= x"0000";
            Ram2(694) <= x"0000";
            Ram2(695) <= x"0000";
            Ram2(696) <= x"0000";
            Ram2(697) <= x"0000";
            Ram2(698) <= x"0000";
            Ram2(699) <= x"0000";
            Ram2(700) <= x"0000";
            Ram2(701) <= x"0000";
            Ram2(702) <= x"0000";
            Ram2(703) <= x"0000";
            Ram2(704) <= x"0000";
            Ram2(705) <= x"0000";
            Ram2(706) <= x"0000";
            Ram2(707) <= x"0000";
            Ram2(708) <= x"0000";
            Ram2(709) <= x"0000";
            Ram2(710) <= x"0000";
            Ram2(711) <= x"0000";
            Ram2(712) <= x"0000";
            Ram2(713) <= x"0000";
            Ram2(714) <= x"0000";
            Ram2(715) <= x"0000";
            Ram2(716) <= x"0000";
            Ram2(717) <= x"0000";
            Ram2(718) <= x"0000";
            Ram2(719) <= x"0000";
            Ram2(720) <= x"0000";
            Ram2(721) <= x"0000";
            Ram2(722) <= x"0000";
            Ram2(723) <= x"0000";
            Ram2(724) <= x"0000";
            Ram2(725) <= x"0000";
            Ram2(726) <= x"0000";
            Ram2(727) <= x"0000";
            Ram2(728) <= x"0000";
            Ram2(729) <= x"0000";
            Ram2(730) <= x"0000";
            Ram2(731) <= x"0000";
            Ram2(732) <= x"0000";
            Ram2(733) <= x"0000";
            Ram2(734) <= x"0000";
            Ram2(735) <= x"0000";
            Ram2(736) <= x"0000";
            Ram2(737) <= x"0000";
            Ram2(738) <= x"0000";
            Ram2(739) <= x"0000";
            Ram2(740) <= x"0000";
            Ram2(741) <= x"0000";
            Ram2(742) <= x"0000";
            Ram2(743) <= x"0000";
            Ram2(744) <= x"0000";
            Ram2(745) <= x"0000";
            Ram2(746) <= x"0000";
            Ram2(747) <= x"0000";
            Ram2(748) <= x"0000";
            Ram2(749) <= x"0000";
            Ram2(750) <= x"0000";
            Ram2(751) <= x"0000";
            Ram2(752) <= x"0000";
            Ram2(753) <= x"0000";
            Ram2(754) <= x"0000";
            Ram2(755) <= x"0000";
            Ram2(756) <= x"0000";
            Ram2(757) <= x"0000";
            Ram2(758) <= x"0000";
            Ram2(759) <= x"0000";
            Ram2(760) <= x"0000";
            Ram2(761) <= x"0000";
            Ram2(762) <= x"0000";
            Ram2(763) <= x"0000";
            Ram2(764) <= x"0000";
            Ram2(765) <= x"0000";
            Ram2(766) <= x"0000";
            Ram2(767) <= x"0000";
            Ram2(768) <= x"0000";
            Ram2(769) <= x"0000";
            Ram2(770) <= x"0000";
            Ram2(771) <= x"0000";
            Ram2(772) <= x"0000";
            Ram2(773) <= x"0000";
            Ram2(774) <= x"0000";
            Ram2(775) <= x"0000";
            Ram2(776) <= x"0000";
            Ram2(777) <= x"0000";
            Ram2(778) <= x"0000";
            Ram2(779) <= x"0000";
            Ram2(780) <= x"0000";
            Ram2(781) <= x"0000";
            Ram2(782) <= x"0000";
            Ram2(783) <= x"0000";
            Ram2(784) <= x"0000";
            Ram2(785) <= x"0000";
            Ram2(786) <= x"0000";
            Ram2(787) <= x"0000";
            Ram2(788) <= x"0000";
            Ram2(789) <= x"0000";
            Ram2(790) <= x"0000";
            Ram2(791) <= x"0000";
            Ram2(792) <= x"0000";
            Ram2(793) <= x"0000";
            Ram2(794) <= x"0000";
            Ram2(795) <= x"0000";
            Ram2(796) <= x"0000";
            Ram2(797) <= x"0000";
            Ram2(798) <= x"0000";
            Ram2(799) <= x"0000";
            Ram2(800) <= x"0000";
            Ram2(801) <= x"0000";
            Ram2(802) <= x"0000";
            Ram2(803) <= x"0000";
            Ram2(804) <= x"0000";
            Ram2(805) <= x"0000";
            Ram2(806) <= x"0000";
            Ram2(807) <= x"0000";
            Ram2(808) <= x"0000";
            Ram2(809) <= x"0000";
            Ram2(810) <= x"0000";
            Ram2(811) <= x"0000";
            Ram2(812) <= x"0000";
            Ram2(813) <= x"0000";
            Ram2(814) <= x"0000";
            Ram2(815) <= x"0000";
            Ram2(816) <= x"0000";
            Ram2(817) <= x"0000";
            Ram2(818) <= x"0000";
            Ram2(819) <= x"0000";
            Ram2(820) <= x"0000";
            Ram2(821) <= x"0000";
            Ram2(822) <= x"0000";
            Ram2(823) <= x"0000";
            Ram2(824) <= x"0000";
            Ram2(825) <= x"0000";
            Ram2(826) <= x"0000";
            Ram2(827) <= x"0000";
            Ram2(828) <= x"0000";
            Ram2(829) <= x"0000";
            Ram2(830) <= x"0000";
            Ram2(831) <= x"0000";
            Ram2(832) <= x"0000";
            Ram2(833) <= x"0000";
            Ram2(834) <= x"0000";
            Ram2(835) <= x"0000";
            Ram2(836) <= x"0000";
            Ram2(837) <= x"0000";
            Ram2(838) <= x"0000";
            Ram2(839) <= x"0000";
            Ram2(840) <= x"0000";
            Ram2(841) <= x"0000";
            Ram2(842) <= x"0000";
            Ram2(843) <= x"0000";
            Ram2(844) <= x"0000";
            Ram2(845) <= x"0000";
            Ram2(846) <= x"0000";
            Ram2(847) <= x"0000";
            Ram2(848) <= x"0000";
            Ram2(849) <= x"0000";
            Ram2(850) <= x"0000";
            Ram2(851) <= x"0000";
            Ram2(852) <= x"0000";
            Ram2(853) <= x"0000";
            Ram2(854) <= x"0000";
            Ram2(855) <= x"0000";
            Ram2(856) <= x"0000";
            Ram2(857) <= x"0000";
            Ram2(858) <= x"0000";
            Ram2(859) <= x"0000";
            Ram2(860) <= x"0000";
            Ram2(861) <= x"0000";
            Ram2(862) <= x"0000";
            Ram2(863) <= x"0000";
            Ram2(864) <= x"0000";
            Ram2(865) <= x"0000";
            Ram2(866) <= x"0000";
            Ram2(867) <= x"0000";
            Ram2(868) <= x"0000";
            Ram2(869) <= x"0000";
            Ram2(870) <= x"0000";
            Ram2(871) <= x"0000";
            Ram2(872) <= x"0000";
            Ram2(873) <= x"0000";
            Ram2(874) <= x"0000";
            Ram2(875) <= x"0000";
            Ram2(876) <= x"0000";
            Ram2(877) <= x"0000";
            Ram2(878) <= x"0000";
            Ram2(879) <= x"0000";
            Ram2(880) <= x"0000";
            Ram2(881) <= x"0000";
            Ram2(882) <= x"0000";
            Ram2(883) <= x"0000";
            Ram2(884) <= x"0000";
            Ram2(885) <= x"0000";
            Ram2(886) <= x"0000";
            Ram2(887) <= x"0000";
            Ram2(888) <= x"0000";
            Ram2(889) <= x"0000";
            Ram2(890) <= x"0000";
            Ram2(891) <= x"0000";
            Ram2(892) <= x"0000";
            Ram2(893) <= x"0000";
            Ram2(894) <= x"0000";
            Ram2(895) <= x"0000";
            Ram2(896) <= x"0000";
            Ram2(897) <= x"0000";
            Ram2(898) <= x"0000";
            Ram2(899) <= x"0000";
            Ram2(900) <= x"0000";
            Ram2(901) <= x"0000";
            Ram2(902) <= x"0000";
            Ram2(903) <= x"0000";
            Ram2(904) <= x"0000";
            Ram2(905) <= x"0000";
            Ram2(906) <= x"0000";
            Ram2(907) <= x"0000";
            Ram2(908) <= x"0000";
            Ram2(909) <= x"0000";
            Ram2(910) <= x"0000";
            Ram2(911) <= x"0000";
            Ram2(912) <= x"0000";
            Ram2(913) <= x"0000";
            Ram2(914) <= x"0000";
            Ram2(915) <= x"0000";
            Ram2(916) <= x"0000";
            Ram2(917) <= x"0000";
            Ram2(918) <= x"0000";
            Ram2(919) <= x"0000";
            Ram2(920) <= x"0000";
            Ram2(921) <= x"0000";
            Ram2(922) <= x"0000";
            Ram2(923) <= x"0000";
            Ram2(924) <= x"0000";
            Ram2(925) <= x"0000";
            Ram2(926) <= x"0000";
            Ram2(927) <= x"0000";
            Ram2(928) <= x"0000";
            Ram2(929) <= x"0000";
            Ram2(930) <= x"0000";
            Ram2(931) <= x"0000";
            Ram2(932) <= x"0000";
            Ram2(933) <= x"0000";
            Ram2(934) <= x"0000";
            Ram2(935) <= x"0000";
            Ram2(936) <= x"0000";
            Ram2(937) <= x"0000";
            Ram2(938) <= x"0000";
            Ram2(939) <= x"0000";
            Ram2(940) <= x"0000";
            Ram2(941) <= x"0000";
            Ram2(942) <= x"0000";
            Ram2(943) <= x"0000";
            Ram2(944) <= x"0000";
            Ram2(945) <= x"0000";
            Ram2(946) <= x"0000";
            Ram2(947) <= x"0000";
            Ram2(948) <= x"0000";
            Ram2(949) <= x"0000";
            Ram2(950) <= x"0000";
            Ram2(951) <= x"0000";
            Ram2(952) <= x"0000";
            Ram2(953) <= x"0000";
            Ram2(954) <= x"0000";
            Ram2(955) <= x"0000";
            Ram2(956) <= x"0000";
            Ram2(957) <= x"0000";
            Ram2(958) <= x"0000";
            Ram2(959) <= x"0000";
            Ram2(960) <= x"0000";
            Ram2(961) <= x"0000";
            Ram2(962) <= x"0000";
            Ram2(963) <= x"0000";
            Ram2(964) <= x"0000";
            Ram2(965) <= x"0000";
            Ram2(966) <= x"0000";
            Ram2(967) <= x"0000";
            Ram2(968) <= x"0000";
            Ram2(969) <= x"0000";
            Ram2(970) <= x"0000";
            Ram2(971) <= x"0000";
            Ram2(972) <= x"0000";
            Ram2(973) <= x"0000";
            Ram2(974) <= x"0000";
            Ram2(975) <= x"0000";
            Ram2(976) <= x"0000";
            Ram2(977) <= x"0000";
            Ram2(978) <= x"0000";
            Ram2(979) <= x"0000";
            Ram2(980) <= x"0000";
            Ram2(981) <= x"0000";
            Ram2(982) <= x"0000";
            Ram2(983) <= x"0000";
            Ram2(984) <= x"0000";
            Ram2(985) <= x"0000";
            Ram2(986) <= x"0000";
            Ram2(987) <= x"0000";
            Ram2(988) <= x"0000";
            Ram2(989) <= x"0000";
            Ram2(990) <= x"0000";
            Ram2(991) <= x"0000";
            Ram2(992) <= x"0000";
            Ram2(993) <= x"0000";
            Ram2(994) <= x"0000";
            Ram2(995) <= x"0000";
            Ram2(996) <= x"0000";
            Ram2(997) <= x"0000";
            Ram2(998) <= x"0000";
            Ram2(999) <= x"0000";
            Ram2(1000) <= x"0000";
            Ram2(1001) <= x"0000";
            Ram2(1002) <= x"0000";
            Ram2(1003) <= x"0000";
            Ram2(1004) <= x"0000";
            Ram2(1005) <= x"0000";
            Ram2(1006) <= x"0000";
            Ram2(1007) <= x"0000";
            Ram2(1008) <= x"0000";
            Ram2(1009) <= x"0000";
            Ram2(1010) <= x"0000";
            Ram2(1011) <= x"0000";
            Ram2(1012) <= x"0000";
            Ram2(1013) <= x"0000";
            Ram2(1014) <= x"0000";
            Ram2(1015) <= x"0000";
            Ram2(1016) <= x"0000";
            Ram2(1017) <= x"0000";
            Ram2(1018) <= x"0000";
            Ram2(1019) <= x"0000";
            Ram2(1020) <= x"0000";
            Ram2(1021) <= x"0000";
            Ram2(1022) <= x"0000";
            Ram2(1023) <= x"0000";
            Ram1(0) <= x"0000";
            Ram1(1) <= x"0000";
            Ram1(2) <= x"0000";
            Ram1(3) <= x"0000";
            Ram1(4) <= x"0000";
            Ram1(5) <= x"0000";
            Ram1(6) <= x"0000";
            Ram1(7) <= x"0000";
            Ram1(8) <= x"0000";
            Ram1(9) <= x"0000";
            Ram1(10) <= x"0000";
            Ram1(11) <= x"0000";
            Ram1(12) <= x"0000";
            Ram1(13) <= x"0000";
            Ram1(14) <= x"0000";
            Ram1(15) <= x"0000";
            Ram1(16) <= x"0000";
            Ram1(17) <= x"0000";
            Ram1(18) <= x"0000";
            Ram1(19) <= x"0000";
            Ram1(20) <= x"0000";
            Ram1(21) <= x"0000";
            Ram1(22) <= x"0000";
            Ram1(23) <= x"0000";
            Ram1(24) <= x"0000";
            Ram1(25) <= x"0000";
            Ram1(26) <= x"0000";
            Ram1(27) <= x"0000";
            Ram1(28) <= x"0000";
            Ram1(29) <= x"0000";
            Ram1(30) <= x"0000";
            Ram1(31) <= x"0000";
            Ram1(32) <= x"0000";
            Ram1(33) <= x"0000";
            Ram1(34) <= x"0000";
            Ram1(35) <= x"0000";
            Ram1(36) <= x"0000";
            Ram1(37) <= x"0000";
            Ram1(38) <= x"0000";
            Ram1(39) <= x"0000";
            Ram1(40) <= x"0000";
            Ram1(41) <= x"0000";
            Ram1(42) <= x"0000";
            Ram1(43) <= x"0000";
            Ram1(44) <= x"0000";
            Ram1(45) <= x"0000";
            Ram1(46) <= x"0000";
            Ram1(47) <= x"0000";
            Ram1(48) <= x"0000";
            Ram1(49) <= x"0000";
            Ram1(50) <= x"0000";
            Ram1(51) <= x"0000";
            Ram1(52) <= x"0000";
            Ram1(53) <= x"0000";
            Ram1(54) <= x"0000";
            Ram1(55) <= x"0000";
            Ram1(56) <= x"0000";
            Ram1(57) <= x"0000";
            Ram1(58) <= x"0000";
            Ram1(59) <= x"0000";
            Ram1(60) <= x"0000";
            Ram1(61) <= x"0000";
            Ram1(62) <= x"0000";
            Ram1(63) <= x"0000";
            Ram1(64) <= x"0000";
            Ram1(65) <= x"0000";
            Ram1(66) <= x"0000";
            Ram1(67) <= x"0000";
            Ram1(68) <= x"0000";
            Ram1(69) <= x"0000";
            Ram1(70) <= x"0000";
            Ram1(71) <= x"0000";
            Ram1(72) <= x"0000";
            Ram1(73) <= x"0000";
            Ram1(74) <= x"0000";
            Ram1(75) <= x"0000";
            Ram1(76) <= x"0000";
            Ram1(77) <= x"0000";
            Ram1(78) <= x"0000";
            Ram1(79) <= x"0000";
            Ram1(80) <= x"0000";
            Ram1(81) <= x"0000";
            Ram1(82) <= x"0000";
            Ram1(83) <= x"0000";
            Ram1(84) <= x"0000";
            Ram1(85) <= x"0000";
            Ram1(86) <= x"0000";
            Ram1(87) <= x"0000";
            Ram1(88) <= x"0000";
            Ram1(89) <= x"0000";
            Ram1(90) <= x"0000";
            Ram1(91) <= x"0000";
            Ram1(92) <= x"0000";
            Ram1(93) <= x"0000";
            Ram1(94) <= x"0000";
            Ram1(95) <= x"0000";
            Ram1(96) <= x"0000";
            Ram1(97) <= x"0000";
            Ram1(98) <= x"0000";
            Ram1(99) <= x"0000";
            Ram1(100) <= x"0000";
            Ram1(101) <= x"0000";
            Ram1(102) <= x"0000";
            Ram1(103) <= x"0000";
            Ram1(104) <= x"0000";
            Ram1(105) <= x"0000";
            Ram1(106) <= x"0000";
            Ram1(107) <= x"0000";
            Ram1(108) <= x"0000";
            Ram1(109) <= x"0000";
            Ram1(110) <= x"0000";
            Ram1(111) <= x"0000";
            Ram1(112) <= x"0000";
            Ram1(113) <= x"0000";
            Ram1(114) <= x"0000";
            Ram1(115) <= x"0000";
            Ram1(116) <= x"0000";
            Ram1(117) <= x"0000";
            Ram1(118) <= x"0000";
            Ram1(119) <= x"0000";
            Ram1(120) <= x"0000";
            Ram1(121) <= x"0000";
            Ram1(122) <= x"0000";
            Ram1(123) <= x"0000";
            Ram1(124) <= x"0000";
            Ram1(125) <= x"0000";
            Ram1(126) <= x"0000";
            Ram1(127) <= x"0000";
            Ram1(128) <= x"0000";
            Ram1(129) <= x"0000";
            Ram1(130) <= x"0000";
            Ram1(131) <= x"0000";
            Ram1(132) <= x"0000";
            Ram1(133) <= x"0000";
            Ram1(134) <= x"0000";
            Ram1(135) <= x"0000";
            Ram1(136) <= x"0000";
            Ram1(137) <= x"0000";
            Ram1(138) <= x"0000";
            Ram1(139) <= x"0000";
            Ram1(140) <= x"0000";
            Ram1(141) <= x"0000";
            Ram1(142) <= x"0000";
            Ram1(143) <= x"0000";
            Ram1(144) <= x"0000";
            Ram1(145) <= x"0000";
            Ram1(146) <= x"0000";
            Ram1(147) <= x"0000";
            Ram1(148) <= x"0000";
            Ram1(149) <= x"0000";
            Ram1(150) <= x"0000";
            Ram1(151) <= x"0000";
            Ram1(152) <= x"0000";
            Ram1(153) <= x"0000";
            Ram1(154) <= x"0000";
            Ram1(155) <= x"0000";
            Ram1(156) <= x"0000";
            Ram1(157) <= x"0000";
            Ram1(158) <= x"0000";
            Ram1(159) <= x"0000";
            Ram1(160) <= x"0000";
            Ram1(161) <= x"0000";
            Ram1(162) <= x"0000";
            Ram1(163) <= x"0000";
            Ram1(164) <= x"0000";
            Ram1(165) <= x"0000";
            Ram1(166) <= x"0000";
            Ram1(167) <= x"0000";
            Ram1(168) <= x"0000";
            Ram1(169) <= x"0000";
            Ram1(170) <= x"0000";
            Ram1(171) <= x"0000";
            Ram1(172) <= x"0000";
            Ram1(173) <= x"0000";
            Ram1(174) <= x"0000";
            Ram1(175) <= x"0000";
            Ram1(176) <= x"0000";
            Ram1(177) <= x"0000";
            Ram1(178) <= x"0000";
            Ram1(179) <= x"0000";
            Ram1(180) <= x"0000";
            Ram1(181) <= x"0000";
            Ram1(182) <= x"0000";
            Ram1(183) <= x"0000";
            Ram1(184) <= x"0000";
            Ram1(185) <= x"0000";
            Ram1(186) <= x"0000";
            Ram1(187) <= x"0000";
            Ram1(188) <= x"0000";
            Ram1(189) <= x"0000";
            Ram1(190) <= x"0000";
            Ram1(191) <= x"0000";
            Ram1(192) <= x"0000";
            Ram1(193) <= x"0000";
            Ram1(194) <= x"0000";
            Ram1(195) <= x"0000";
            Ram1(196) <= x"0000";
            Ram1(197) <= x"0000";
            Ram1(198) <= x"0000";
            Ram1(199) <= x"0000";
            Ram1(200) <= x"0000";
            Ram1(201) <= x"0000";
            Ram1(202) <= x"0000";
            Ram1(203) <= x"0000";
            Ram1(204) <= x"0000";
            Ram1(205) <= x"0000";
            Ram1(206) <= x"0000";
            Ram1(207) <= x"0000";
            Ram1(208) <= x"0000";
            Ram1(209) <= x"0000";
            Ram1(210) <= x"0000";
            Ram1(211) <= x"0000";
            Ram1(212) <= x"0000";
            Ram1(213) <= x"0000";
            Ram1(214) <= x"0000";
            Ram1(215) <= x"0000";
            Ram1(216) <= x"0000";
            Ram1(217) <= x"0000";
            Ram1(218) <= x"0000";
            Ram1(219) <= x"0000";
            Ram1(220) <= x"0000";
            Ram1(221) <= x"0000";
            Ram1(222) <= x"0000";
            Ram1(223) <= x"0000";
            Ram1(224) <= x"0000";
            Ram1(225) <= x"0000";
            Ram1(226) <= x"0000";
            Ram1(227) <= x"0000";
            Ram1(228) <= x"0000";
            Ram1(229) <= x"0000";
            Ram1(230) <= x"0000";
            Ram1(231) <= x"0000";
            Ram1(232) <= x"0000";
            Ram1(233) <= x"0000";
            Ram1(234) <= x"0000";
            Ram1(235) <= x"0000";
            Ram1(236) <= x"0000";
            Ram1(237) <= x"0000";
            Ram1(238) <= x"0000";
            Ram1(239) <= x"0000";
            Ram1(240) <= x"0000";
            Ram1(241) <= x"0000";
            Ram1(242) <= x"0000";
            Ram1(243) <= x"0000";
            Ram1(244) <= x"0000";
            Ram1(245) <= x"0000";
            Ram1(246) <= x"0000";
            Ram1(247) <= x"0000";
            Ram1(248) <= x"0000";
            Ram1(249) <= x"0000";
            Ram1(250) <= x"0000";
            Ram1(251) <= x"0000";
            Ram1(252) <= x"0000";
            Ram1(253) <= x"0000";
            Ram1(254) <= x"0000";
            Ram1(255) <= x"0000";
            Ram1(256) <= x"0000";
            Ram1(257) <= x"0000";
            Ram1(258) <= x"0000";
            Ram1(259) <= x"0000";
            Ram1(260) <= x"0000";
            Ram1(261) <= x"0000";
            Ram1(262) <= x"0000";
            Ram1(263) <= x"0000";
            Ram1(264) <= x"0000";
            Ram1(265) <= x"0000";
            Ram1(266) <= x"0000";
            Ram1(267) <= x"0000";
            Ram1(268) <= x"0000";
            Ram1(269) <= x"0000";
            Ram1(270) <= x"0000";
            Ram1(271) <= x"0000";
            Ram1(272) <= x"0000";
            Ram1(273) <= x"0000";
            Ram1(274) <= x"0000";
            Ram1(275) <= x"0000";
            Ram1(276) <= x"0000";
            Ram1(277) <= x"0000";
            Ram1(278) <= x"0000";
            Ram1(279) <= x"0000";
            Ram1(280) <= x"0000";
            Ram1(281) <= x"0000";
            Ram1(282) <= x"0000";
            Ram1(283) <= x"0000";
            Ram1(284) <= x"0000";
            Ram1(285) <= x"0000";
            Ram1(286) <= x"0000";
            Ram1(287) <= x"0000";
            Ram1(288) <= x"0000";
            Ram1(289) <= x"0000";
            Ram1(290) <= x"0000";
            Ram1(291) <= x"0000";
            Ram1(292) <= x"0000";
            Ram1(293) <= x"0000";
            Ram1(294) <= x"0000";
            Ram1(295) <= x"0000";
            Ram1(296) <= x"0000";
            Ram1(297) <= x"0000";
            Ram1(298) <= x"0000";
            Ram1(299) <= x"0000";
            Ram1(300) <= x"0000";
            Ram1(301) <= x"0000";
            Ram1(302) <= x"0000";
            Ram1(303) <= x"0000";
            Ram1(304) <= x"0000";
            Ram1(305) <= x"0000";
            Ram1(306) <= x"0000";
            Ram1(307) <= x"0000";
            Ram1(308) <= x"0000";
            Ram1(309) <= x"0000";
            Ram1(310) <= x"0000";
            Ram1(311) <= x"0000";
            Ram1(312) <= x"0000";
            Ram1(313) <= x"0000";
            Ram1(314) <= x"0000";
            Ram1(315) <= x"0000";
            Ram1(316) <= x"0000";
            Ram1(317) <= x"0000";
            Ram1(318) <= x"0000";
            Ram1(319) <= x"0000";
            Ram1(320) <= x"0000";
            Ram1(321) <= x"0000";
            Ram1(322) <= x"0000";
            Ram1(323) <= x"0000";
            Ram1(324) <= x"0000";
            Ram1(325) <= x"0000";
            Ram1(326) <= x"0000";
            Ram1(327) <= x"0000";
            Ram1(328) <= x"0000";
            Ram1(329) <= x"0000";
            Ram1(330) <= x"0000";
            Ram1(331) <= x"0000";
            Ram1(332) <= x"0000";
            Ram1(333) <= x"0000";
            Ram1(334) <= x"0000";
            Ram1(335) <= x"0000";
            Ram1(336) <= x"0000";
            Ram1(337) <= x"0000";
            Ram1(338) <= x"0000";
            Ram1(339) <= x"0000";
            Ram1(340) <= x"0000";
            Ram1(341) <= x"0000";
            Ram1(342) <= x"0000";
            Ram1(343) <= x"0000";
            Ram1(344) <= x"0000";
            Ram1(345) <= x"0000";
            Ram1(346) <= x"0000";
            Ram1(347) <= x"0000";
            Ram1(348) <= x"0000";
            Ram1(349) <= x"0000";
            Ram1(350) <= x"0000";
            Ram1(351) <= x"0000";
            Ram1(352) <= x"0000";
            Ram1(353) <= x"0000";
            Ram1(354) <= x"0000";
            Ram1(355) <= x"0000";
            Ram1(356) <= x"0000";
            Ram1(357) <= x"0000";
            Ram1(358) <= x"0000";
            Ram1(359) <= x"0000";
            Ram1(360) <= x"0000";
            Ram1(361) <= x"0000";
            Ram1(362) <= x"0000";
            Ram1(363) <= x"0000";
            Ram1(364) <= x"0000";
            Ram1(365) <= x"0000";
            Ram1(366) <= x"0000";
            Ram1(367) <= x"0000";
            Ram1(368) <= x"0000";
            Ram1(369) <= x"0000";
            Ram1(370) <= x"0000";
            Ram1(371) <= x"0000";
            Ram1(372) <= x"0000";
            Ram1(373) <= x"0000";
            Ram1(374) <= x"0000";
            Ram1(375) <= x"0000";
            Ram1(376) <= x"0000";
            Ram1(377) <= x"0000";
            Ram1(378) <= x"0000";
            Ram1(379) <= x"0000";
            Ram1(380) <= x"0000";
            Ram1(381) <= x"0000";
            Ram1(382) <= x"0000";
            Ram1(383) <= x"0000";
            Ram1(384) <= x"0000";
            Ram1(385) <= x"0000";
            Ram1(386) <= x"0000";
            Ram1(387) <= x"0000";
            Ram1(388) <= x"0000";
            Ram1(389) <= x"0000";
            Ram1(390) <= x"0000";
            Ram1(391) <= x"0000";
            Ram1(392) <= x"0000";
            Ram1(393) <= x"0000";
            Ram1(394) <= x"0000";
            Ram1(395) <= x"0000";
            Ram1(396) <= x"0000";
            Ram1(397) <= x"0000";
            Ram1(398) <= x"0000";
            Ram1(399) <= x"0000";
            Ram1(400) <= x"0000";
            Ram1(401) <= x"0000";
            Ram1(402) <= x"0000";
            Ram1(403) <= x"0000";
            Ram1(404) <= x"0000";
            Ram1(405) <= x"0000";
            Ram1(406) <= x"0000";
            Ram1(407) <= x"0000";
            Ram1(408) <= x"0000";
            Ram1(409) <= x"0000";
            Ram1(410) <= x"0000";
            Ram1(411) <= x"0000";
            Ram1(412) <= x"0000";
            Ram1(413) <= x"0000";
            Ram1(414) <= x"0000";
            Ram1(415) <= x"0000";
            Ram1(416) <= x"0000";
            Ram1(417) <= x"0000";
            Ram1(418) <= x"0000";
            Ram1(419) <= x"0000";
            Ram1(420) <= x"0000";
            Ram1(421) <= x"0000";
            Ram1(422) <= x"0000";
            Ram1(423) <= x"0000";
            Ram1(424) <= x"0000";
            Ram1(425) <= x"0000";
            Ram1(426) <= x"0000";
            Ram1(427) <= x"0000";
            Ram1(428) <= x"0000";
            Ram1(429) <= x"0000";
            Ram1(430) <= x"0000";
            Ram1(431) <= x"0000";
            Ram1(432) <= x"0000";
            Ram1(433) <= x"0000";
            Ram1(434) <= x"0000";
            Ram1(435) <= x"0000";
            Ram1(436) <= x"0000";
            Ram1(437) <= x"0000";
            Ram1(438) <= x"0000";
            Ram1(439) <= x"0000";
            Ram1(440) <= x"0000";
            Ram1(441) <= x"0000";
            Ram1(442) <= x"0000";
            Ram1(443) <= x"0000";
            Ram1(444) <= x"0000";
            Ram1(445) <= x"0000";
            Ram1(446) <= x"0000";
            Ram1(447) <= x"0000";
            Ram1(448) <= x"0000";
            Ram1(449) <= x"0000";
            Ram1(450) <= x"0000";
            Ram1(451) <= x"0000";
            Ram1(452) <= x"0000";
            Ram1(453) <= x"0000";
            Ram1(454) <= x"0000";
            Ram1(455) <= x"0000";
            Ram1(456) <= x"0000";
            Ram1(457) <= x"0000";
            Ram1(458) <= x"0000";
            Ram1(459) <= x"0000";
            Ram1(460) <= x"0000";
            Ram1(461) <= x"0000";
            Ram1(462) <= x"0000";
            Ram1(463) <= x"0000";
            Ram1(464) <= x"0000";
            Ram1(465) <= x"0000";
            Ram1(466) <= x"0000";
            Ram1(467) <= x"0000";
            Ram1(468) <= x"0000";
            Ram1(469) <= x"0000";
            Ram1(470) <= x"0000";
            Ram1(471) <= x"0000";
            Ram1(472) <= x"0000";
            Ram1(473) <= x"0000";
            Ram1(474) <= x"0000";
            Ram1(475) <= x"0000";
            Ram1(476) <= x"0000";
            Ram1(477) <= x"0000";
            Ram1(478) <= x"0000";
            Ram1(479) <= x"0000";
            Ram1(480) <= x"0000";
            Ram1(481) <= x"0000";
            Ram1(482) <= x"0000";
            Ram1(483) <= x"0000";
            Ram1(484) <= x"0000";
            Ram1(485) <= x"0000";
            Ram1(486) <= x"0000";
            Ram1(487) <= x"0000";
            Ram1(488) <= x"0000";
            Ram1(489) <= x"0000";
            Ram1(490) <= x"0000";
            Ram1(491) <= x"0000";
            Ram1(492) <= x"0000";
            Ram1(493) <= x"0000";
            Ram1(494) <= x"0000";
            Ram1(495) <= x"0000";
            Ram1(496) <= x"0000";
            Ram1(497) <= x"0000";
            Ram1(498) <= x"0000";
            Ram1(499) <= x"0000";
            Ram1(500) <= x"0000";
            Ram1(501) <= x"0000";
            Ram1(502) <= x"0000";
            Ram1(503) <= x"0000";
            Ram1(504) <= x"0000";
            Ram1(505) <= x"0000";
            Ram1(506) <= x"0000";
            Ram1(507) <= x"0000";
            Ram1(508) <= x"0000";
            Ram1(509) <= x"0000";
            Ram1(510) <= x"0000";
            Ram1(511) <= x"0000";
            Ram1(512) <= x"0000";
            Ram1(513) <= x"0000";
            Ram1(514) <= x"0000";
            Ram1(515) <= x"0000";
            Ram1(516) <= x"0000";
            Ram1(517) <= x"0000";
            Ram1(518) <= x"0000";
            Ram1(519) <= x"0000";
            Ram1(520) <= x"0000";
            Ram1(521) <= x"0000";
            Ram1(522) <= x"0000";
            Ram1(523) <= x"0000";
            Ram1(524) <= x"0000";
            Ram1(525) <= x"0000";
            Ram1(526) <= x"0000";
            Ram1(527) <= x"0000";
            Ram1(528) <= x"0000";
            Ram1(529) <= x"0000";
            Ram1(530) <= x"0000";
            Ram1(531) <= x"0000";
            Ram1(532) <= x"0000";
            Ram1(533) <= x"0000";
            Ram1(534) <= x"0000";
            Ram1(535) <= x"0000";
            Ram1(536) <= x"0000";
            Ram1(537) <= x"0000";
            Ram1(538) <= x"0000";
            Ram1(539) <= x"0000";
            Ram1(540) <= x"0000";
            Ram1(541) <= x"0000";
            Ram1(542) <= x"0000";
            Ram1(543) <= x"0000";
            Ram1(544) <= x"0000";
            Ram1(545) <= x"0000";
            Ram1(546) <= x"0000";
            Ram1(547) <= x"0000";
            Ram1(548) <= x"0000";
            Ram1(549) <= x"0000";
            Ram1(550) <= x"0000";
            Ram1(551) <= x"0000";
            Ram1(552) <= x"0000";
            Ram1(553) <= x"0000";
            Ram1(554) <= x"0000";
            Ram1(555) <= x"0000";
            Ram1(556) <= x"0000";
            Ram1(557) <= x"0000";
            Ram1(558) <= x"0000";
            Ram1(559) <= x"0000";
            Ram1(560) <= x"0000";
            Ram1(561) <= x"0000";
            Ram1(562) <= x"0000";
            Ram1(563) <= x"0000";
            Ram1(564) <= x"0000";
            Ram1(565) <= x"0000";
            Ram1(566) <= x"0000";
            Ram1(567) <= x"0000";
            Ram1(568) <= x"0000";
            Ram1(569) <= x"0000";
            Ram1(570) <= x"0000";
            Ram1(571) <= x"0000";
            Ram1(572) <= x"0000";
            Ram1(573) <= x"0000";
            Ram1(574) <= x"0000";
            Ram1(575) <= x"0000";
            Ram1(576) <= x"0000";
            Ram1(577) <= x"0000";
            Ram1(578) <= x"0000";
            Ram1(579) <= x"0000";
            Ram1(580) <= x"0000";
            Ram1(581) <= x"0000";
            Ram1(582) <= x"0000";
            Ram1(583) <= x"0000";
            Ram1(584) <= x"0000";
            Ram1(585) <= x"0000";
            Ram1(586) <= x"0000";
            Ram1(587) <= x"0000";
            Ram1(588) <= x"0000";
            Ram1(589) <= x"0000";
            Ram1(590) <= x"0000";
            Ram1(591) <= x"0000";
            Ram1(592) <= x"0000";
            Ram1(593) <= x"0000";
            Ram1(594) <= x"0000";
            Ram1(595) <= x"0000";
            Ram1(596) <= x"0000";
            Ram1(597) <= x"0000";
            Ram1(598) <= x"0000";
            Ram1(599) <= x"0000";
            Ram1(600) <= x"0000";
            Ram1(601) <= x"0000";
            Ram1(602) <= x"0000";
            Ram1(603) <= x"0000";
            Ram1(604) <= x"0000";
            Ram1(605) <= x"0000";
            Ram1(606) <= x"0000";
            Ram1(607) <= x"0000";
            Ram1(608) <= x"0000";
            Ram1(609) <= x"0000";
            Ram1(610) <= x"0000";
            Ram1(611) <= x"0000";
            Ram1(612) <= x"0000";
            Ram1(613) <= x"0000";
            Ram1(614) <= x"0000";
            Ram1(615) <= x"0000";
            Ram1(616) <= x"0000";
            Ram1(617) <= x"0000";
            Ram1(618) <= x"0000";
            Ram1(619) <= x"0000";
            Ram1(620) <= x"0000";
            Ram1(621) <= x"0000";
            Ram1(622) <= x"0000";
            Ram1(623) <= x"0000";
            Ram1(624) <= x"0000";
            Ram1(625) <= x"0000";
            Ram1(626) <= x"0000";
            Ram1(627) <= x"0000";
            Ram1(628) <= x"0000";
            Ram1(629) <= x"0000";
            Ram1(630) <= x"0000";
            Ram1(631) <= x"0000";
            Ram1(632) <= x"0000";
            Ram1(633) <= x"0000";
            Ram1(634) <= x"0000";
            Ram1(635) <= x"0000";
            Ram1(636) <= x"0000";
            Ram1(637) <= x"0000";
            Ram1(638) <= x"0000";
            Ram1(639) <= x"0000";
            Ram1(640) <= x"0000";
            Ram1(641) <= x"0000";
            Ram1(642) <= x"0000";
            Ram1(643) <= x"0000";
            Ram1(644) <= x"0000";
            Ram1(645) <= x"0000";
            Ram1(646) <= x"0000";
            Ram1(647) <= x"0000";
            Ram1(648) <= x"0000";
            Ram1(649) <= x"0000";
            Ram1(650) <= x"0000";
            Ram1(651) <= x"0000";
            Ram1(652) <= x"0000";
            Ram1(653) <= x"0000";
            Ram1(654) <= x"0000";
            Ram1(655) <= x"0000";
            Ram1(656) <= x"0000";
            Ram1(657) <= x"0000";
            Ram1(658) <= x"0000";
            Ram1(659) <= x"0000";
            Ram1(660) <= x"0000";
            Ram1(661) <= x"0000";
            Ram1(662) <= x"0000";
            Ram1(663) <= x"0000";
            Ram1(664) <= x"0000";
            Ram1(665) <= x"0000";
            Ram1(666) <= x"0000";
            Ram1(667) <= x"0000";
            Ram1(668) <= x"0000";
            Ram1(669) <= x"0000";
            Ram1(670) <= x"0000";
            Ram1(671) <= x"0000";
            Ram1(672) <= x"0000";
            Ram1(673) <= x"0000";
            Ram1(674) <= x"0000";
            Ram1(675) <= x"0000";
            Ram1(676) <= x"0000";
            Ram1(677) <= x"0000";
            Ram1(678) <= x"0000";
            Ram1(679) <= x"0000";
            Ram1(680) <= x"0000";
            Ram1(681) <= x"0000";
            Ram1(682) <= x"0000";
            Ram1(683) <= x"0000";
            Ram1(684) <= x"0000";
            Ram1(685) <= x"0000";
            Ram1(686) <= x"0000";
            Ram1(687) <= x"0000";
            Ram1(688) <= x"0000";
            Ram1(689) <= x"0000";
            Ram1(690) <= x"0000";
            Ram1(691) <= x"0000";
            Ram1(692) <= x"0000";
            Ram1(693) <= x"0000";
            Ram1(694) <= x"0000";
            Ram1(695) <= x"0000";
            Ram1(696) <= x"0000";
            Ram1(697) <= x"0000";
            Ram1(698) <= x"0000";
            Ram1(699) <= x"0000";
            Ram1(700) <= x"0000";
            Ram1(701) <= x"0000";
            Ram1(702) <= x"0000";
            Ram1(703) <= x"0000";
            Ram1(704) <= x"0000";
            Ram1(705) <= x"0000";
            Ram1(706) <= x"0000";
            Ram1(707) <= x"0000";
            Ram1(708) <= x"0000";
            Ram1(709) <= x"0000";
            Ram1(710) <= x"0000";
            Ram1(711) <= x"0000";
            Ram1(712) <= x"0000";
            Ram1(713) <= x"0000";
            Ram1(714) <= x"0000";
            Ram1(715) <= x"0000";
            Ram1(716) <= x"0000";
            Ram1(717) <= x"0000";
            Ram1(718) <= x"0000";
            Ram1(719) <= x"0000";
            Ram1(720) <= x"0000";
            Ram1(721) <= x"0000";
            Ram1(722) <= x"0000";
            Ram1(723) <= x"0000";
            Ram1(724) <= x"0000";
            Ram1(725) <= x"0000";
            Ram1(726) <= x"0000";
            Ram1(727) <= x"0000";
            Ram1(728) <= x"0000";
            Ram1(729) <= x"0000";
            Ram1(730) <= x"0000";
            Ram1(731) <= x"0000";
            Ram1(732) <= x"0000";
            Ram1(733) <= x"0000";
            Ram1(734) <= x"0000";
            Ram1(735) <= x"0000";
            Ram1(736) <= x"0000";
            Ram1(737) <= x"0000";
            Ram1(738) <= x"0000";
            Ram1(739) <= x"0000";
            Ram1(740) <= x"0000";
            Ram1(741) <= x"0000";
            Ram1(742) <= x"0000";
            Ram1(743) <= x"0000";
            Ram1(744) <= x"0000";
            Ram1(745) <= x"0000";
            Ram1(746) <= x"0000";
            Ram1(747) <= x"0000";
            Ram1(748) <= x"0000";
            Ram1(749) <= x"0000";
            Ram1(750) <= x"0000";
            Ram1(751) <= x"0000";
            Ram1(752) <= x"0000";
            Ram1(753) <= x"0000";
            Ram1(754) <= x"0000";
            Ram1(755) <= x"0000";
            Ram1(756) <= x"0000";
            Ram1(757) <= x"0000";
            Ram1(758) <= x"0000";
            Ram1(759) <= x"0000";
            Ram1(760) <= x"0000";
            Ram1(761) <= x"0000";
            Ram1(762) <= x"0000";
            Ram1(763) <= x"0000";
            Ram1(764) <= x"0000";
            Ram1(765) <= x"0000";
            Ram1(766) <= x"0000";
            Ram1(767) <= x"0000";
            Ram1(768) <= x"0000";
            Ram1(769) <= x"0000";
            Ram1(770) <= x"0000";
            Ram1(771) <= x"0000";
            Ram1(772) <= x"0000";
            Ram1(773) <= x"0000";
            Ram1(774) <= x"0000";
            Ram1(775) <= x"0000";
            Ram1(776) <= x"0000";
            Ram1(777) <= x"0000";
            Ram1(778) <= x"0000";
            Ram1(779) <= x"0000";
            Ram1(780) <= x"0000";
            Ram1(781) <= x"0000";
            Ram1(782) <= x"0000";
            Ram1(783) <= x"0000";
            Ram1(784) <= x"0000";
            Ram1(785) <= x"0000";
            Ram1(786) <= x"0000";
            Ram1(787) <= x"0000";
            Ram1(788) <= x"0000";
            Ram1(789) <= x"0000";
            Ram1(790) <= x"0000";
            Ram1(791) <= x"0000";
            Ram1(792) <= x"0000";
            Ram1(793) <= x"0000";
            Ram1(794) <= x"0000";
            Ram1(795) <= x"0000";
            Ram1(796) <= x"0000";
            Ram1(797) <= x"0000";
            Ram1(798) <= x"0000";
            Ram1(799) <= x"0000";
            Ram1(800) <= x"0000";
            Ram1(801) <= x"0000";
            Ram1(802) <= x"0000";
            Ram1(803) <= x"0000";
            Ram1(804) <= x"0000";
            Ram1(805) <= x"0000";
            Ram1(806) <= x"0000";
            Ram1(807) <= x"0000";
            Ram1(808) <= x"0000";
            Ram1(809) <= x"0000";
            Ram1(810) <= x"0000";
            Ram1(811) <= x"0000";
            Ram1(812) <= x"0000";
            Ram1(813) <= x"0000";
            Ram1(814) <= x"0000";
            Ram1(815) <= x"0000";
            Ram1(816) <= x"0000";
            Ram1(817) <= x"0000";
            Ram1(818) <= x"0000";
            Ram1(819) <= x"0000";
            Ram1(820) <= x"0000";
            Ram1(821) <= x"0000";
            Ram1(822) <= x"0000";
            Ram1(823) <= x"0000";
            Ram1(824) <= x"0000";
            Ram1(825) <= x"0000";
            Ram1(826) <= x"0000";
            Ram1(827) <= x"0000";
            Ram1(828) <= x"0000";
            Ram1(829) <= x"0000";
            Ram1(830) <= x"0000";
            Ram1(831) <= x"0000";
            Ram1(832) <= x"0000";
            Ram1(833) <= x"0000";
            Ram1(834) <= x"0000";
            Ram1(835) <= x"0000";
            Ram1(836) <= x"0000";
            Ram1(837) <= x"0000";
            Ram1(838) <= x"0000";
            Ram1(839) <= x"0000";
            Ram1(840) <= x"0000";
            Ram1(841) <= x"0000";
            Ram1(842) <= x"0000";
            Ram1(843) <= x"0000";
            Ram1(844) <= x"0000";
            Ram1(845) <= x"0000";
            Ram1(846) <= x"0000";
            Ram1(847) <= x"0000";
            Ram1(848) <= x"0000";
            Ram1(849) <= x"0000";
            Ram1(850) <= x"0000";
            Ram1(851) <= x"0000";
            Ram1(852) <= x"0000";
            Ram1(853) <= x"0000";
            Ram1(854) <= x"0000";
            Ram1(855) <= x"0000";
            Ram1(856) <= x"0000";
            Ram1(857) <= x"0000";
            Ram1(858) <= x"0000";
            Ram1(859) <= x"0000";
            Ram1(860) <= x"0000";
            Ram1(861) <= x"0000";
            Ram1(862) <= x"0000";
            Ram1(863) <= x"0000";
            Ram1(864) <= x"0000";
            Ram1(865) <= x"0000";
            Ram1(866) <= x"0000";
            Ram1(867) <= x"0000";
            Ram1(868) <= x"0000";
            Ram1(869) <= x"0000";
            Ram1(870) <= x"0000";
            Ram1(871) <= x"0000";
            Ram1(872) <= x"0000";
            Ram1(873) <= x"0000";
            Ram1(874) <= x"0000";
            Ram1(875) <= x"0000";
            Ram1(876) <= x"0000";
            Ram1(877) <= x"0000";
            Ram1(878) <= x"0000";
            Ram1(879) <= x"0000";
            Ram1(880) <= x"0000";
            Ram1(881) <= x"0000";
            Ram1(882) <= x"0000";
            Ram1(883) <= x"0000";
            Ram1(884) <= x"0000";
            Ram1(885) <= x"0000";
            Ram1(886) <= x"0000";
            Ram1(887) <= x"0000";
            Ram1(888) <= x"0000";
            Ram1(889) <= x"0000";
            Ram1(890) <= x"0000";
            Ram1(891) <= x"0000";
            Ram1(892) <= x"0000";
            Ram1(893) <= x"0000";
            Ram1(894) <= x"0000";
            Ram1(895) <= x"0000";
            Ram1(896) <= x"0000";
            Ram1(897) <= x"0000";
            Ram1(898) <= x"0000";
            Ram1(899) <= x"0000";
            Ram1(900) <= x"0000";
            Ram1(901) <= x"0000";
            Ram1(902) <= x"0000";
            Ram1(903) <= x"0000";
            Ram1(904) <= x"0000";
            Ram1(905) <= x"0000";
            Ram1(906) <= x"0000";
            Ram1(907) <= x"0000";
            Ram1(908) <= x"0000";
            Ram1(909) <= x"0000";
            Ram1(910) <= x"0000";
            Ram1(911) <= x"0000";
            Ram1(912) <= x"0000";
            Ram1(913) <= x"0000";
            Ram1(914) <= x"0000";
            Ram1(915) <= x"0000";
            Ram1(916) <= x"0000";
            Ram1(917) <= x"0000";
            Ram1(918) <= x"0000";
            Ram1(919) <= x"0000";
            Ram1(920) <= x"0000";
            Ram1(921) <= x"0000";
            Ram1(922) <= x"0000";
            Ram1(923) <= x"0000";
            Ram1(924) <= x"0000";
            Ram1(925) <= x"0000";
            Ram1(926) <= x"0000";
            Ram1(927) <= x"0000";
            Ram1(928) <= x"0000";
            Ram1(929) <= x"0000";
            Ram1(930) <= x"0000";
            Ram1(931) <= x"0000";
            Ram1(932) <= x"0000";
            Ram1(933) <= x"0000";
            Ram1(934) <= x"0000";
            Ram1(935) <= x"0000";
            Ram1(936) <= x"0000";
            Ram1(937) <= x"0000";
            Ram1(938) <= x"0000";
            Ram1(939) <= x"0000";
            Ram1(940) <= x"0000";
            Ram1(941) <= x"0000";
            Ram1(942) <= x"0000";
            Ram1(943) <= x"0000";
            Ram1(944) <= x"0000";
            Ram1(945) <= x"0000";
            Ram1(946) <= x"0000";
            Ram1(947) <= x"0000";
            Ram1(948) <= x"0000";
            Ram1(949) <= x"0000";
            Ram1(950) <= x"0000";
            Ram1(951) <= x"0000";
            Ram1(952) <= x"0000";
            Ram1(953) <= x"0000";
            Ram1(954) <= x"0000";
            Ram1(955) <= x"0000";
            Ram1(956) <= x"0000";
            Ram1(957) <= x"0000";
            Ram1(958) <= x"0000";
            Ram1(959) <= x"0000";
            Ram1(960) <= x"0000";
            Ram1(961) <= x"0000";
            Ram1(962) <= x"0000";
            Ram1(963) <= x"0000";
            Ram1(964) <= x"0000";
            Ram1(965) <= x"0000";
            Ram1(966) <= x"0000";
            Ram1(967) <= x"0000";
            Ram1(968) <= x"0000";
            Ram1(969) <= x"0000";
            Ram1(970) <= x"0000";
            Ram1(971) <= x"0000";
            Ram1(972) <= x"0000";
            Ram1(973) <= x"0000";
            Ram1(974) <= x"0000";
            Ram1(975) <= x"0000";
            Ram1(976) <= x"0000";
            Ram1(977) <= x"0000";
            Ram1(978) <= x"0000";
            Ram1(979) <= x"0000";
            Ram1(980) <= x"0000";
            Ram1(981) <= x"0000";
            Ram1(982) <= x"0000";
            Ram1(983) <= x"0000";
            Ram1(984) <= x"0000";
            Ram1(985) <= x"0000";
            Ram1(986) <= x"0000";
            Ram1(987) <= x"0000";
            Ram1(988) <= x"0000";
            Ram1(989) <= x"0000";
            Ram1(990) <= x"0000";
            Ram1(991) <= x"0000";
            Ram1(992) <= x"0000";
            Ram1(993) <= x"0000";
            Ram1(994) <= x"0000";
            Ram1(995) <= x"0000";
            Ram1(996) <= x"0000";
            Ram1(997) <= x"0000";
            Ram1(998) <= x"0000";
            Ram1(999) <= x"0000";
            Ram1(1000) <= x"0000";
            Ram1(1001) <= x"0000";
            Ram1(1002) <= x"0000";
            Ram1(1003) <= x"0000";
            Ram1(1004) <= x"0000";
            Ram1(1005) <= x"0000";
            Ram1(1006) <= x"0000";
            Ram1(1007) <= x"0000";
            Ram1(1008) <= x"0000";
            Ram1(1009) <= x"0000";
            Ram1(1010) <= x"0000";
            Ram1(1011) <= x"0000";
            Ram1(1012) <= x"0000";
            Ram1(1013) <= x"0000";
            Ram1(1014) <= x"0000";
            Ram1(1015) <= x"0000";
            Ram1(1016) <= x"0000";
            Ram1(1017) <= x"0000";
            Ram1(1018) <= x"0000";
            Ram1(1019) <= x"0000";
            Ram1(1020) <= x"0000";
            Ram1(1021) <= x"0000";
            Ram1(1022) <= x"0000";
            Ram1(1023) <= x"0000";
		elsif (clk_scan'event and clk_scan = '1' and startedCache = '1') then
			if (triggercache /= (LFlag & SFlag & Address & DataS & InstructionAddress)) then
				triggerCache <= LFlag & SFlag & Address & DataS & InstructionAddress;
				if (((LFlag or SFlag) = '1') and Address < x"8000") then
					if (LFlag = '1') then
						Result <= Ram2(conv_integer(Address(9 downto 0)));
						Result_L <= Ram2(conv_integer(Address(9 downto 0)));
						Result_L_pointer <= '1';
					else
						Ram2(conv_integer(Address(9 downto 0))) <= DataS;
						Result <= (others => '0');
						Result_L <= (others => '0');
						Result_L_pointer <= '0';
					end if;
					InstructionResult <= (others => '0');
				else
					InstructionResult <= Ram2(conv_integer(InstructionAddress(9 downto 0)));
					if (LFlag = '1') then
						Result <= Ram1(conv_integer(Address(9 downto 0)));
						Result_L <= Ram1(conv_integer(Address(9 downto 0)));
						Result_L_pointer <= '1';
					elsif (SFlag = '1') then
						Ram1(conv_integer(Address(9 downto 0))) <= DataS;
						Result <= (others => '0');
						Result_L <= (others => '0');
						Result_L_pointer <= '1';
					else
						Result <= Address;
						Result_L <= Address;
						Result_L_pointer <= '0';
					end if;
				end if;
			end if;
		end if;
	end process;
end bhv;