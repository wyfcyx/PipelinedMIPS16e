library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity main is
	port(
		clk : in std_logic;
		output : out std_logic_vector(1 downto 0)
	);
end main;

architecture bhv of main is

begin

end bhv;

